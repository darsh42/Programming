module chip8 (clock, reset);

   input clock;
   input reset;



endmodule // chip8

module 1NNN (PC, CIR)
   inout [16:0] PC;
   input [16:0] CIR;


endmodule // 1NNN
